module tbGlobal_tb;
  //global testbench code
endmodule
